library verilog;
use verilog.vl_types.all;
entity ULA8bits_vlg_vec_tst is
end ULA8bits_vlg_vec_tst;
